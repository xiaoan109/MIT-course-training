import Types::*;
import ProcTypes::*;
import CacheTypes::*;
import MemTypes::*;
import Fifo::*;
import Vector::*;

module mkParentProtocolProcessor(MessageFifo#(n) r2m, MessageFifo#(n) m2r, WideMem mem, Empty ifc);
    // TODO: implement the parent protocol processor
endmodule

